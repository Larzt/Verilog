module ul4 (output wire[3:0] Out, input wire[3:0] A, input wire[3:0] B, input wire [1:0] S);
endmodule